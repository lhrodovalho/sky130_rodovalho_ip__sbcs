* NGSPICE file created from bjt.ext - technology: sky130A

.subckt sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 Emitter Collector Base m=1
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
.ends

.subckt bjt x
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
+ VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
.ends

