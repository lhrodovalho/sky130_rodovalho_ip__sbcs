magic
tech sky130A
timestamp 1717055877
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1715908107
transform 1 0 0 0 1 0
box 0 0 670 670
<< end >>
