* expanding   symbol:  sbcs0.sym # of pins=7
* sym_path: /home/rodovalho/git/sky130_rodovalho_ip__sbcs/xschem/sbcs0.sym
* sch_path: /home/rodovalho/git/sky130_rodovalho_ip__sbcs/xschem/sbcs0.sch
.subckt sbcs0  isource  isink  en  enb  avdd  avss  vsub
*.iopin isink
*.iopin isource
*.ipin enb
*.ipin en
*.iopin avss
*.iopin avdd
*.iopin vsub
xslice[1] isource isink en enb avdd avss vsub bpa0 bpa bpb x y bn0 bn z sbcs0_slice
xslice[0] isource isink en enb avdd avss vsub bpa0 bpa bpb x y bn0 bn z sbcs0_slice
.ends


* expanding   symbol:  sbcs0_slice.sym # of pins=15
* sym_path: /home/rodovalho/git/sky130_rodovalho_ip__sbcs/xschem/sbcs0_slice.sym
* sch_path: /home/rodovalho/git/sky130_rodovalho_ip__sbcs/xschem/sbcs0_slice.sch
.subckt sbcs0_slice  isource  isink  en  enb  avdd  avss  vsub  bpa0  bpa  bpb  x  y  bn0  bn  z
*.iopin isink
*.iopin isource
*.ipin enb
*.ipin en
*.iopin avss
*.iopin avdd
*.iopin bpb
*.iopin bpa
*.iopin bn
*.iopin x
*.iopin y
*.iopin bn0
*.iopin bpa0
*.iopin vsub
*.iopin z
x1c bn0 bn0 y avss n1_1
x2d bpa0 bn0 avss avss n1_2
x3d bpa bn avss avss n1_2
x1b bn0 bpb w1a avdd p1_2
x1a w1a bpa avdd avdd p1_2
x2b bpa0 bpb w2a avdd p1_2
x2a w2a bpa0 avdd avdd p1_2
x3b bpa bpb w3a avdd p1_2
x3a w3a bpa0 avdd avdd p1_2
x5d bn bn avss avss n1_2
x5b bn_ bpb w5a avdd p1_2
x5a w5a bpa avdd avdd p1_2
x6d bpb bn avss avss n2_1
x6a_ bpb bpb avdd avdd p1_4
x9b isource bpb w9a avdd p2_1
x9a w9a bpa avdd avdd p2_1
x8d z bn avss avss n1_1
x7c w7b z bn avss n1_1
x7b avdd en w7b avss n1_1
x4d_ bn enb avss avss n1_1
x5c bn_ en bn avss n1_1
x4a bpa en avdd avdd p1_2
x7a avdd z avdd avdd p1_2
x8a z en avdd avdd p1_1
x9d isink bn avss avss n2_1
XR1 avss y avss sky130_fd_pr__res_xhigh_po W=1 L=5.7 mult=1 m=1
.ends


* expanding   symbol:  n1_1.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130_rodovalho_ip__sbcs/xschem/n1_1.sym
* sch_path: /home/rodovalho/git/sky130_rodovalho_ip__sbcs/xschem/n1_1.sch
.subckt n1_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XMD[3] D G X[3] B sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMD[2] D G X[2] B sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMD[1] D G X[1] B sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMD[0] D G X[0] B sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMS[3] X[3] G S B sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMS[2] X[2] G S B sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMS[1] X[1] G S B sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMS[0] X[0] G S B sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  n1_2.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130_rodovalho_ip__sbcs/xschem/n1_2.sym
* sch_path: /home/rodovalho/git/sky130_rodovalho_ip__sbcs/xschem/n1_2.sch
.subckt n1_2  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xd D G X B n1_1
xs X G S B n1_1
.ends


* expanding   symbol:  p1_2.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130_rodovalho_ip__sbcs/xschem/p1_2.sym
* sch_path: /home/rodovalho/git/sky130_rodovalho_ip__sbcs/xschem/p1_2.sch
.subckt p1_2  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xs X G S B p1_1
xd D G X B p1_1
.ends


* expanding   symbol:  n2_1.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130_rodovalho_ip__sbcs/xschem/n2_1.sym
* sch_path: /home/rodovalho/git/sky130_rodovalho_ip__sbcs/xschem/n2_1.sch
.subckt n2_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xr D G S B n1_1
xl D G S B n1_1
.ends


* expanding   symbol:  p1_4.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130_rodovalho_ip__sbcs/xschem/p1_4.sym
* sch_path: /home/rodovalho/git/sky130_rodovalho_ip__sbcs/xschem/p1_4.sch
.subckt p1_4  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xs X G S B p1_2
xd D G X B p1_2
.ends


* expanding   symbol:  p2_1.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130_rodovalho_ip__sbcs/xschem/p2_1.sym
* sch_path: /home/rodovalho/git/sky130_rodovalho_ip__sbcs/xschem/p2_1.sch
.subckt p2_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xl D G S B p1_1
xr D G S B p1_1
.ends


* expanding   symbol:  p1_1.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130_rodovalho_ip__sbcs/xschem/p1_1.sym
* sch_path: /home/rodovalho/git/sky130_rodovalho_ip__sbcs/xschem/p1_1.sch
.subckt p1_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM0[7] D G S B sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=5.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM0[6] D G S B sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=5.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM0[5] D G S B sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=5.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM0[4] D G S B sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=5.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM0[3] D G S B sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=5.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM0[2] D G S B sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=5.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM0[1] D G S B sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=5.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM0[0] D G S B sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=5.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends
